library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

package synchronizer_pkg is

    type coefficients is array(natural range <>) of signed(15 downto 0);

end package synchronizer_pkg;
